`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:28:16 04/13/2019 
// Design Name: 
// Module Name:    writer 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module writer(
    input Clock,
    input [7:0] Data,
    input [7:0] Address,
    output SDA,
    output SCL,
    output Busy
    );


endmodule
